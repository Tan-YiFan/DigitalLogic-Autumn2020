`ifndef __LAB6_SVH
`define __LAB6_SVH



`endif

module decoder2_4 (
    input logic [1:0] in,
    output logic [3:0] out,
    input logic en
);
    
endmodule

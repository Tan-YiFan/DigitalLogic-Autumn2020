module ans (
    input logic [3:0]in,
    output logic [6:0]out
);
    always_comb begin
        unique case(in)
            
            default: begin
                
            end
        endcase
    end
    
endmodule

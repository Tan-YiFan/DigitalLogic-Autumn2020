module top (
    input logic clk, resetn,
    output logic LED16_G, LED16_R, LED17_G
);
endmodule

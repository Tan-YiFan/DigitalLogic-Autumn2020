module lab6 (
    
);

endmodule

module lab4 (
    input logic [3:0]in,
    output logic [6:0]out_use138, out_use151
);
    seg_138 seg_138_inst(.in, .out(out_use138));
    seg_151 seg_151_inst(.in, .out(out_use151));
endmodule

module seg_138 (
    input logic [3:0]in,
    output logic [6:0]out
);
    // TODO: add logic here
    // NOTE: "always_comb" are not allowed here. You should use mod_74LS138 instants and logic gates(assign) here

endmodule

module mod_74LS138 (
    // TODO: add ports here

);
    // TODO: add logic here
    // NOTE: No syntax limitation

endmodule

module seg_151 (
    input logic [3:0]in,
    output logic [6:0]out
);
    // TODO: add logic here
    // NOTE: "always_comb" are not allowed here. You should use mod_74LS151 instants and logic gates(assign) here

endmodule

module mod_74LS151 (
    // TODO: add ports here
    
);
    // TODO: add logic here
    // NOTE: No syntax limitation

endmodule
module sim (
    
);
endmodule

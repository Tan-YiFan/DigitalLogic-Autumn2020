module lab2 (
    input logic [31:0]instr,
    output logic [7:0]aluout
);
    // TODO: add signal declaration here

    decoder myDecoder(
        // TODO: add ports here
    );

    alu myALU(
        // TODO: add ports here
    );

endmodule

module decoder (
    // TODO: add port declaration here

);
    // TODO: add logic here

endmodule

module alu (
    // TODO: add port declaration here
);
    // TODO: add logic here

endmodule

module sim (
    
);
    
    decoder4_16 sim1();
    decoder5_32 sim2();
    encoder16_4 sim3();
    priority_encoder16_4 sim4();
endmodule

`ifndef __DECODER_SVH
`define __DECODER_SVH



`endif

module priority_encoder4_2 (
    input logic [3:0] in,
    output logic [1:0] out
);
    
endmodule

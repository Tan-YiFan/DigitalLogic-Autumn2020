module lab7 (
    input logic clk,
    // ...

);

endmodule

module sim (
    
);

endmodule

module top (
    input logic clk, resetn,
    output logic LED16_G, LED_16_R, LED17_G, LED17_R,
    output logic [6:0]A2G,
    output logic [7:0]AN
);

endmodule
